package router_test_pkg;
     import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "router_wr_xtn.sv"
    `include "source_config.sv"
    `include "dest_config.sv"
    `include "env_config.sv"
    `include "source_driver.sv"
    `include "source_monitor.sv"
    `include "source_sequencer.sv"
    `include "source_agent.sv"
    `include "source_agent_top.sv"
    `include "source_sequence.sv"
    
    `include "router_rd_xtn.sv"
    `include "dest_driver.sv"
    `include "dest_monitor.sv"
    `include "dest_sequencer.sv"
    `include "dst_agent.sv"
    `include "dest_agt_top.sv"
    `include "dest_sequences.sv" 
       
    `include "virtual_seqr.sv"
    `include "virtual_seqs.sv"
     
    `include "router_scoreboard.sv"
    `include "router_env.sv"
    `include "router_test.sv"
endpackage
